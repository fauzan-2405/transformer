// linear_projection.sv
// Used to do linear projection of course (duh)
import linear_proj_pkg::*;

module linear_pojection #(
    parameter XXX = YY
) (
    input logic xxx,
    output logic yyy
);
    // Bismillah

endmodule