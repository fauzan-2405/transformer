// multi_matmul.v
// Used to wrap multi matmul module

module multi_matmul #(
    parameter siuuuu = 2
) (
    input clk,
    input rst_n
);
    localparam euyyyy = 3;

endmodule