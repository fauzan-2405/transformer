// softmax_lut.v
// Used to store LUT values 
// The input ranges from -8 to +8
// Output is in Q16.16 fixed-point format: [S][15 INT][16 FRAC]

module softmax_lut #(
    parameter WIDTH = 16,
    parameter FRAC_WIDTH = 8,
    parameter INT_WIDTH = 8
) (
    input  wire signed [INT_WIDTH-1:0] in,      // Range: -8 to +8
    output reg  [WIDTH*2-1:0] e_i_val          
);
    always @(*) begin
        case (in)
            -8: e_i_val = 32'b0000000000000000_0000000000010110; // 22       ≈ 0.00033546
            -7: e_i_val = 32'b0000000000000000_0000000001011110; // 94       ≈ 0.00183156
            -6: e_i_val = 32'b0000000000000000_0000000011111011; // 507      ≈ 0.00773619
            -5: e_i_val = 32'b0000000000000000_0000001010111000; // 1368     ≈ 0.02087402
            -4: e_i_val = 32'b0000000000000000_0000011011011100; // 3548     ≈ 0.05407715
            -3: e_i_val = 32'b0000000000000000_0001001111111001; // 5113     ≈ 0.07803345
            -2: e_i_val = 32'b0000000000000000_0010001011011110; // 8798     ≈ 0.13429260
            -1: e_i_val = 32'b0000000000000000_0101111100001101; // 24397    ≈ 0.37243652
             0: e_i_val = 32'b0000000000000001_0000000000000000; // 65536    = 1.0
             1: e_i_val = 32'b0000000000000010_1011100001010001; // 178145   ≈ 2.71828
             2: e_i_val = 32'b0000000000000111_0110001110011011; // 483099   ≈ 7.38906
             3: e_i_val = 32'b0000000000010100_0001001011110010; // 1318050  ≈ 20.0855
             4: e_i_val = 32'b0000000000110110_1000100111111000; // 3575528  ≈ 54.5982
             5: e_i_val = 32'b0000000010010100_1111100110111000; // 9732096  ≈ 148.413
             6: e_i_val = 32'b0000001011001010_1111011110011000; // 26424184 ≈ 403.429
             7: e_i_val = 32'b0000010001001110_1011101111101011; // 71839819 ≈ 1096.63
             8: e_i_val = 32'b0000101110101111_1111000000000111; // 195105927 ≈ 2980.96
            default: e_i_val = 32'b0000000000000000_0000000000000000; // default = 0
        endcase
    end
endmodule
