// matmul_linear_proj.v
// Used to do linear projection for Q, K, and V

module matmul_linear_proj #(
    parameter siuuuu = 2
) (
    input clk,
    input rst_n
);
    localparam euyyyy = 3;

endmodule