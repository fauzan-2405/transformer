// top_linear_projection.sv
// Top module for linear_projection (keys + matmul modules) + controller + input BRAM
import linear_proj_pkg::*;

module top_linear_projection #(
    parameter XXXX = yy
) (
    input logic clk,
    output logic xxx
);

endmodule