// top_self_attention_head.sv
// This is the top module for self_attention_head + self_attention_ctrl

module top_self_attention_head #(
    parameter XXX = YYY
) (
    input logic clk, rst_n,

    output logic xxx
);
    
endmodule