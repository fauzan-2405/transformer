// bridge_buffer_ctrl.sv
// Used to control bridge_buffer
// Basically utilizing the linear_proj_ctrl.sv but tweaks some of the settings

module bridge_buffer_ctrl #(
    parameter XXX = YYY,
    parameter XXX = YYY,
) (
    input logic clk, rst_n,
    output logic xxx
);
    

endmodule