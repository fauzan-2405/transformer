// linear_projection.v
// Used to do linear projection for Q, K, and V

module linear_projection #(
    parameter siuuuu = 2
) (
    input clk,
    input rst_n
);
    localparam euyyyy = 3;
    
endmodule