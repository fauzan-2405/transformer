// This package contains parameters used in self attention head 

package self_attention_pkg;
    
endpackage