// multwrap_wbram.sv
// This used to wrap multi_matmul_wrapper.sv + its corresponding BRAM