module blockmatmul
  (
    
  )
